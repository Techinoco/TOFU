
module CMA ( CLK, RST_N, CBANK, RUN, EXWE, EXRE, EXWD, EXROMUL, EXA, DBGSEL, 
        EXRD, DBGDAT, DONE, CLK_FOR_ARRAY );
  input [24:0] EXWD;
  input [19:0] EXROMUL;
  input [11:0] EXA;
  input [2:0] DBGSEL;
  output [24:0] EXRD;
  output [3:0] DBGDAT;
  input CLK, RST_N, CBANK, RUN, EXWE, EXRE, CLK_FOR_ARRAY;
  output DONE;

  wire   [299:0] TOPEARRAY;
  wire   [299:0] FPEARRAY;
  wire   [383:0] CONF_ALU;
  wire   [287:0] CONF_SEL_A;
  wire   [287:0] CONF_SEL_B;
  wire   [959:0] CONF_SE;
  wire   [135:0] CONST_DATA_A;
  wire   [135:0] CONST_DATA_B;

  // mc mc1 ( .CLK(CLK), .RST_N(RST_N), .CBANK(CBANK), .RUN(RUN), .TOPEARRAY(
  //       TOPEARRAY), .FPEARRAY(FPEARRAY), .CONF_ALU(CONF_ALU), .CONF_SEL_A(
  //       CONF_SEL_A), .CONF_SEL_B(CONF_SEL_B), .CONF_SE(CONF_SE), 
  //       .CONST_DATA_A(CONST_DATA_A), .CONST_DATA_B(CONST_DATA_B), .DONE(DONE), 
  //       .EXWE(EXWE), .EXRE(EXRE), .EXWD(EXWD), .EXRD(EXRD), .EXROMUL(EXROMUL), 
  //       .EXA(EXA), .DBGSEL(DBGSEL), .DBGDAT(DBGDAT) );
mc mc1(
    .CLK (CLK), .RST_N(RST_N), .CBANK(CBANK), .RUN(RUN),
    .TOPEARRAY     (TOPEARRAY),
    .FPEARRAY      (FPEARRAY),// SWOPED D3
    .CONF_ALU      (CONF_ALU),
    .CONF_SEL_A    (CONF_SEL_A),
    .CONF_SEL_B    (CONF_SEL_B),
    .CONF_SE       (CONF_SE),
    .CONST_DATA_A  (CONST_DATA_A),
    .CONST_DATA_B  (CONST_DATA_B),
    .DONE          (DONE),
    .EXWE          (EXWE), 
    .EXRE          (EXRE),
    .EXWD          (EXWD),
    .EXRD          (EXRD),
    .EXROMUL       (EXROMUL),
    .EXA           (EXA),
    .DBGSEL        (DBGSEL),
    .DBGDAT        (DBGDAT)
);
PE_ARRAY PE_ARRAY1 (
    .CLK           (CLK_FOR_ARRAY),
    .RST_N         (RST_N),
    .CONF_ALU      (CONF_ALU),
    .CONF_SEL_A    (CONF_SEL_A),
    .CONF_SEL_B    (CONF_SEL_B),
    .CONF_SE       (CONF_SE),
    .IN_SOUTH      (TOPEARRAY),
    .IN_CONST_A    (CONST_DATA_A),
    .IN_CONST_B    (CONST_DATA_B),
    .OUT_SOUTH     (FPEARRAY)
);
  // PE_ARRAY PE_ARRAY1 ( .CLK(CLK), .RST_N(RST_N), .CONF_ALU(CONF_ALU), .CONF_SEL_A(CONF_SEL_A), .CONF_SEL_B(CONF_SEL_B), .CONF_SE(CONF_SE), .IN_SOUTH(TOPEARRAY), 
  //       .IN_CONST_A(CONST_DATA_A), .IN_CONST_B(CONST_DATA_B), .OUT_SOUTH(
  //       FPEARRAY) );
endmodule

module CMA_TOP (EXWD,EXROMUL,EXA,DBGSEL,EXRD,DBGDAT,CLK,RST_N,CBANK,RUN,EXWE,EXRE,CLK_FOR_ARRAY,DONE);
	wire [24:0] EXWD_int;
	input [24:0] EXWD;
	wire [19:0] EXROMUL_int;
	input [19:0] EXROMUL;
	wire [11:0] EXA_int;
	input [11:0] EXA;
	wire [2:0] DBGSEL_int;
	input [2:0] DBGSEL;
	wire [24:0] EXRD_int;
	output [24:0] EXRD;
	wire [3:0] DBGDAT_int;
	output [3:0] DBGDAT;
	input CLK;
	wire CLK_int;
	input RST_N;
	wire RST_N_int;
	input CBANK;
	wire CBANK_int;
	input RUN;
	wire RUN_int;
	input EXWE;
	wire EXWE_int;
	input EXRE;
	wire EXRE_int;
	input CLK_FOR_ARRAY;
	wire CLK_FOR_ARRAY_int;
	output DONE;
	wire DONE_int;
	LE8HIOT3B02BZ_IN U0_0 (.PAD(EXWD[0]),.CIN(EXWD_int[0]));
	LE8HIOT3B02BZ_IN U0_1 (.PAD(EXWD[1]),.CIN(EXWD_int[1]));
	LE8HIOT3B02BZ_IN U0_2 (.PAD(EXWD[2]),.CIN(EXWD_int[2]));
	LE8HIOT3B02BZ_IN U0_3 (.PAD(EXWD[3]),.CIN(EXWD_int[3]));
	LE8HIOT3B02BZ_IN U0_4 (.PAD(EXWD[4]),.CIN(EXWD_int[4]));
	LE8HIOT3B02BZ_IN U0_5 (.PAD(EXWD[5]),.CIN(EXWD_int[5]));
	LE8HIOT3B02BZ_IN U0_6 (.PAD(EXWD[6]),.CIN(EXWD_int[6]));
	LE8HIOT3B02BZ_IN U0_7 (.PAD(EXWD[7]),.CIN(EXWD_int[7]));
	LE8HIOT3B02BZ_IN U0_8 (.PAD(EXWD[8]),.CIN(EXWD_int[8]));
	LE8HIOT3B02BZ_IN U0_9 (.PAD(EXWD[9]),.CIN(EXWD_int[9]));
	LE8HIOT3B02BZ_IN U0_10 (.PAD(EXWD[10]),.CIN(EXWD_int[10]));
	LE8HIOT3B02BZ_IN U0_11 (.PAD(EXWD[11]),.CIN(EXWD_int[11]));
	LE8HIOT3B02BZ_IN U0_12 (.PAD(EXWD[12]),.CIN(EXWD_int[12]));
	LE8HIOT3B02BZ_IN U0_13 (.PAD(EXWD[13]),.CIN(EXWD_int[13]));
	LE8HIOT3B02BZ_IN U0_14 (.PAD(EXWD[14]),.CIN(EXWD_int[14]));
	LE8HIOT3B02BZ_IN U0_15 (.PAD(EXWD[15]),.CIN(EXWD_int[15]));
	LE8HIOT3B02BZ_IN U0_16 (.PAD(EXWD[16]),.CIN(EXWD_int[16]));
	LE8HIOT3B02BZ_IN U0_17 (.PAD(EXWD[17]),.CIN(EXWD_int[17]));
	LE8HIOT3B02BZ_IN U0_18 (.PAD(EXWD[18]),.CIN(EXWD_int[18]));
	LE8HIOT3B02BZ_IN U0_19 (.PAD(EXWD[19]),.CIN(EXWD_int[19]));
	LE8HIOT3B02BZ_IN U0_20 (.PAD(EXWD[20]),.CIN(EXWD_int[20]));
	LE8HIOT3B02BZ_IN U0_21 (.PAD(EXWD[21]),.CIN(EXWD_int[21]));
	LE8HIOT3B02BZ_IN U0_22 (.PAD(EXWD[22]),.CIN(EXWD_int[22]));
	LE8HIOT3B02BZ_IN U0_23 (.PAD(EXWD[23]),.CIN(EXWD_int[23]));
	LE8HIOT3B02BZ_IN U0_24 (.PAD(EXWD[24]),.CIN(EXWD_int[24]));
	LE8HIOT3B02BZ_IN U1_0 (.PAD(EXROMUL[0]),.CIN(EXROMUL_int[0]));
	LE8HIOT3B02BZ_IN U1_1 (.PAD(EXROMUL[1]),.CIN(EXROMUL_int[1]));
	LE8HIOT3B02BZ_IN U1_2 (.PAD(EXROMUL[2]),.CIN(EXROMUL_int[2]));
	LE8HIOT3B02BZ_IN U1_3 (.PAD(EXROMUL[3]),.CIN(EXROMUL_int[3]));
	LE8HIOT3B02BZ_IN U1_4 (.PAD(EXROMUL[4]),.CIN(EXROMUL_int[4]));
	LE8HIOT3B02BZ_IN U1_5 (.PAD(EXROMUL[5]),.CIN(EXROMUL_int[5]));
	LE8HIOT3B02BZ_IN U1_6 (.PAD(EXROMUL[6]),.CIN(EXROMUL_int[6]));
	LE8HIOT3B02BZ_IN U1_7 (.PAD(EXROMUL[7]),.CIN(EXROMUL_int[7]));
	LE8HIOT3B02BZ_IN U1_8 (.PAD(EXROMUL[8]),.CIN(EXROMUL_int[8]));
	LE8HIOT3B02BZ_IN U1_9 (.PAD(EXROMUL[9]),.CIN(EXROMUL_int[9]));
	LE8HIOT3B02BZ_IN U1_10 (.PAD(EXROMUL[10]),.CIN(EXROMUL_int[10]));
	LE8HIOT3B02BZ_IN U1_11 (.PAD(EXROMUL[11]),.CIN(EXROMUL_int[11]));
	LE8HIOT3B02BZ_IN U1_12 (.PAD(EXROMUL[12]),.CIN(EXROMUL_int[12]));
	LE8HIOT3B02BZ_IN U1_13 (.PAD(EXROMUL[13]),.CIN(EXROMUL_int[13]));
	LE8HIOT3B02BZ_IN U1_14 (.PAD(EXROMUL[14]),.CIN(EXROMUL_int[14]));
	LE8HIOT3B02BZ_IN U1_15 (.PAD(EXROMUL[15]),.CIN(EXROMUL_int[15]));
	LE8HIOT3B02BZ_IN U1_16 (.PAD(EXROMUL[16]),.CIN(EXROMUL_int[16]));
	LE8HIOT3B02BZ_IN U1_17 (.PAD(EXROMUL[17]),.CIN(EXROMUL_int[17]));
	LE8HIOT3B02BZ_IN U1_18 (.PAD(EXROMUL[18]),.CIN(EXROMUL_int[18]));
	LE8HIOT3B02BZ_IN U1_19 (.PAD(EXROMUL[19]),.CIN(EXROMUL_int[19]));
	LE8HIOT3B02BZ_IN U2_0 (.PAD(EXA[0]),.CIN(EXA_int[0]));
	LE8HIOT3B02BZ_IN U2_1 (.PAD(EXA[1]),.CIN(EXA_int[1]));
	LE8HIOT3B02BZ_IN U2_2 (.PAD(EXA[2]),.CIN(EXA_int[2]));
	LE8HIOT3B02BZ_IN U2_3 (.PAD(EXA[3]),.CIN(EXA_int[3]));
	LE8HIOT3B02BZ_IN U2_4 (.PAD(EXA[4]),.CIN(EXA_int[4]));
	LE8HIOT3B02BZ_IN U2_5 (.PAD(EXA[5]),.CIN(EXA_int[5]));
	LE8HIOT3B02BZ_IN U2_6 (.PAD(EXA[6]),.CIN(EXA_int[6]));
	LE8HIOT3B02BZ_IN U2_7 (.PAD(EXA[7]),.CIN(EXA_int[7]));
	LE8HIOT3B02BZ_IN U2_8 (.PAD(EXA[8]),.CIN(EXA_int[8]));
	LE8HIOT3B02BZ_IN U2_9 (.PAD(EXA[9]),.CIN(EXA_int[9]));
	LE8HIOT3B02BZ_IN U2_10 (.PAD(EXA[10]),.CIN(EXA_int[10]));
	LE8HIOT3B02BZ_IN U2_11 (.PAD(EXA[11]),.CIN(EXA_int[11]));
	LE8HIOT3B02BZ_IN U3_0 (.PAD(DBGSEL[0]),.CIN(DBGSEL_int[0]));
	LE8HIOT3B02BZ_IN U3_1 (.PAD(DBGSEL[1]),.CIN(DBGSEL_int[1]));
	LE8HIOT3B02BZ_IN U3_2 (.PAD(DBGSEL[2]),.CIN(DBGSEL_int[2]));
	LE8HIOT3B02BZ_OUT U4_0 (.PAD(EXRD[0]),.I(EXRD_int[0]));
	LE8HIOT3B02BZ_OUT U4_1 (.PAD(EXRD[1]),.I(EXRD_int[1]));
	LE8HIOT3B02BZ_OUT U4_2 (.PAD(EXRD[2]),.I(EXRD_int[2]));
	LE8HIOT3B02BZ_OUT U4_3 (.PAD(EXRD[3]),.I(EXRD_int[3]));
	LE8HIOT3B02BZ_OUT U4_4 (.PAD(EXRD[4]),.I(EXRD_int[4]));
	LE8HIOT3B02BZ_OUT U4_5 (.PAD(EXRD[5]),.I(EXRD_int[5]));
	LE8HIOT3B02BZ_OUT U4_6 (.PAD(EXRD[6]),.I(EXRD_int[6]));
	LE8HIOT3B02BZ_OUT U4_7 (.PAD(EXRD[7]),.I(EXRD_int[7]));
	LE8HIOT3B02BZ_OUT U4_8 (.PAD(EXRD[8]),.I(EXRD_int[8]));
	LE8HIOT3B02BZ_OUT U4_9 (.PAD(EXRD[9]),.I(EXRD_int[9]));
	LE8HIOT3B02BZ_OUT U4_10 (.PAD(EXRD[10]),.I(EXRD_int[10]));
	LE8HIOT3B02BZ_OUT U4_11 (.PAD(EXRD[11]),.I(EXRD_int[11]));
	LE8HIOT3B02BZ_OUT U4_12 (.PAD(EXRD[12]),.I(EXRD_int[12]));
	LE8HIOT3B02BZ_OUT U4_13 (.PAD(EXRD[13]),.I(EXRD_int[13]));
	LE8HIOT3B02BZ_OUT U4_14 (.PAD(EXRD[14]),.I(EXRD_int[14]));
	LE8HIOT3B02BZ_OUT U4_15 (.PAD(EXRD[15]),.I(EXRD_int[15]));
	LE8HIOT3B02BZ_OUT U4_16 (.PAD(EXRD[16]),.I(EXRD_int[16]));
	LE8HIOT3B02BZ_OUT U4_17 (.PAD(EXRD[17]),.I(EXRD_int[17]));
	LE8HIOT3B02BZ_OUT U4_18 (.PAD(EXRD[18]),.I(EXRD_int[18]));
	LE8HIOT3B02BZ_OUT U4_19 (.PAD(EXRD[19]),.I(EXRD_int[19]));
	LE8HIOT3B02BZ_OUT U4_20 (.PAD(EXRD[20]),.I(EXRD_int[20]));
	LE8HIOT3B02BZ_OUT U4_21 (.PAD(EXRD[21]),.I(EXRD_int[21]));
	LE8HIOT3B02BZ_OUT U4_22 (.PAD(EXRD[22]),.I(EXRD_int[22]));
	LE8HIOT3B02BZ_OUT U4_23 (.PAD(EXRD[23]),.I(EXRD_int[23]));
	LE8HIOT3B02BZ_OUT U4_24 (.PAD(EXRD[24]),.I(EXRD_int[24]));
	LE8HIOT3B02BZ_OUT U5_0 (.PAD(DBGDAT[0]),.I(DBGDAT_int[0]));
	LE8HIOT3B02BZ_OUT U5_1 (.PAD(DBGDAT[1]),.I(DBGDAT_int[1]));
	LE8HIOT3B02BZ_OUT U5_2 (.PAD(DBGDAT[2]),.I(DBGDAT_int[2]));
	LE8HIOT3B02BZ_OUT U5_3 (.PAD(DBGDAT[3]),.I(DBGDAT_int[3]));
	LE8HIOT3B02BZ_IN U6 (.PAD(CLK),.CIN(CLK_int));
	LE8HIOT3B02BZ_IN U7 (.PAD(RST_N),.CIN(RST_N_int));
	LE8HIOT3B02BZ_IN U8 (.PAD(CBANK),.CIN(CBANK_int));
	LE8HIOT3B02BZ_IN U9 (.PAD(RUN),.CIN(RUN_int));
	LE8HIOT3B02BZ_IN U10 (.PAD(EXWE),.CIN(EXWE_int));
	LE8HIOT3B02BZ_IN U11 (.PAD(EXRE),.CIN(EXRE_int));
	LE8HIOT3B02BZ_IN U12 (.PAD(CLK_FOR_ARRAY),.CIN(CLK_FOR_ARRAY_int));
	LE8HIOT3B02BZ_OUT U13 (.PAD(DONE),.I(DONE_int));
	CMA I0 (
 		.EXWD(EXWD_int),
 		.EXROMUL(EXROMUL_int),
 		.EXA(EXA_int),
 		.DBGSEL(DBGSEL_int),
 		.EXRD(EXRD_int),
 		.DBGDAT(DBGDAT_int),
 		.CLK(CLK_int),
 		.RST_N(RST_N_int),
 		.CBANK(CBANK_int),
 		.RUN(RUN_int),
 		.EXWE(EXWE_int),
 		.EXRE(EXRE_int),
 		.CLK_FOR_ARRAY(CLK_FOR_ARRAY_int),
 		.DONE(DONE_int));
endmodule
